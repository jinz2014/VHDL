type mem_data_md is array ( 0 to 7, 0 to 3) of std_logic;

constant rom : mem_data_md :=
( 
  ('0', '0', '0', '0'),
  ('0', '0', '0', '1'),
  ('0', '0', '1', '0'),
  ('0', '1', '1', '1'),
  ('0', '1', '0', '0'),
  ('0', '1', '1', '1'),
  ('0', '1', '1', '0'),
  ('0', '1', '1', '1')
);


x := rom(3,3);
